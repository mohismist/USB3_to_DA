library verilog;
use verilog.vl_types.all;
entity sig_pll_altpll is
    port(
        clk             : out    vl_logic_vector(4 downto 0);
        inclk           : in     vl_logic_vector(1 downto 0);
        locked          : out    vl_logic
    );
end sig_pll_altpll;
